LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Test_Alarm IS
	PORT (CLOCK_50: IN STD_LOGIC;
			SW: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			HEX0, HEX1, HEX2: OUT  STD_LOGIC_VECTOR(6 DOWNTO 0));
END Test_Alarm;

ARCHITECTURE BEHAVIOUR OF Test_Alarm IS
Signal clock: STD_LOGIC;
BEGIN

Pre_scale: work.PreScale port map (CLOCK_50, clock);
Test: work.Alarm port map (clock, SW(0), HEX0, HEX1, HEX2);

END BEHAVIOUR;